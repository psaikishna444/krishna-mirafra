class axi_r_driver extends uvm_driver#(axi_transaction);

`uvm_component_utils(axi_r_driver)

//virtual axi_if.RDRV rdvif;
virtual axi_if vif;


axi_transaction rtrans;

int num_sent1;

//constructor//////////

function new(string name="axi_r_driver",uvm_component parent);
super.new(name,parent);
endfunction

function void build_phase(uvm_phase phase);
super.build_phase(phase);
if(!uvm_config_db#(virtual axi_if)::get(this,"","vif",vif))
`uvm_fatal("NO_VIF",{"virtual interface must be set for:",get_full_name(),".vif"});
rtrans=axi_transaction::type_id::create("rtrans",this);
endfunction
///////////////////START OF SIMULATION//////////////////

function void start_of_simulation_phase(uvm_phase phase );
		`uvm_info(get_type_name(),{"start of simulation for ",get_full_name()},UVM_LOW)
	endfunction



//////////////////RUN PHASE/////////////////////////



task run_phase(uvm_phase phase);
 forever
   begin
      repeat(5) @(vif.r_drv_cb);
         if(!vif.r_drv_cb.rst)
           begin      
       		`uvm_info(get_type_name(),"RESET observed",UVM_LOW)
                 vif.r_drv_cb.arvalid <= 0;   
                 vif.r_drv_cb.araddr <= 'bx;   
                 vif.r_drv_cb.arprot <= 0;   
                 vif.r_drv_cb.rready <= 0;
		            end  
         else
          begin

              seq_item_port.get_next_item(rtrans);  
                          vif.r_drv_cb.arvalid <= rtrans.arvalid;  
			//  vif.r_drv_cb.arvalid <= 1'b1;      
		    //repeat (1) @ (vif.r_drv_cb);
                      if(vif.r_drv_cb.arready && vif.r_drv_cb.arvalid) 
                         begin
			 vif.r_drv_cb.araddr <= rtrans.araddr;
    			 vif.r_drv_cb.arprot <= rtrans.arprot;
         vif.r_drv_cb.rready <= rtrans.rready;
	  //vif.r_drv_cb.rready <= 1'b1;	
		num_sent1++;
                         end
		seq_item_port.item_done();

          end
  end			
 endtask  
      

/*
task run_phase (uvm_phase phase);
forever 
begin
repeat(5)@(vif.r_drv_cb);
		if (!vif.r_drv_cb.rst)
	begin
	`uvm_info(get_type_name(),"RESET observed",UVM_LOW)
		vif.r_drv_cb.rdata<=32'hZZZ;
		vif.r_drv_cb.arready<=1'b0;
		vif.r_drv_cb.awready<=1'b0;
		vif.r_drv_cb.wready<=1'b0;
		vif.r_drv_cb.bvalid<=1'b0;
		vif.r_drv_cb.bresp<=1'b0;
		vif.r_drv_cb.araddr<=32'hxx;
		vif.r_drv_cb.arprot<=3'b000;
		vif.r_drv_cb.rvalid<=1'b0;
		vif.r_drv_cb.rresp<=1'b0;
	end
	else

	begin
	seq_item_port.get_next_item(rtrans);
			@(vif.r_drv_cb);

	///////////////////write address channel//////////////

	vif.r_drv_cb.awready<=1'b1;
		@(vif.r_drv_cb);
		wait(vif.r_drv_cb.awvalid);
			@(vif.r_drv_cb);
			vif.r_drv_cb.awready<=1'b0;
			vif.r_drv_cb.awaddr<=rtrans.awaddr;
			vif.r_drv_cb.awprot<=rtrans.awprot;

	//////////////write data //////////////////
	@(vif.r_drv_cb);
		vif.r_drv_cb.wready<=1'b1;
		@(vif.r_drv_cb);
		wait(vif.r_drv_cb.wvalid);
		@(vif.r_drv_cb);
		vif.r_drv_cb.wready<=1'b0;

		vif.r_drv_cb.wdata<=rtrans.wdata;
		vif.r_drv_cb.wstrb<=rtrans.wstrb;

//////////////////////write response/////////////////

	@(vif.r_drv_cb);

		vif.r_drv_cb.bvalid<=1'b1;
		wait(vif.r_drv_cb.bready);
		vif.r_drv_cb.bresp<=1'b1;

	@(vif.r_drv_cb);
	
		vif.r_drv_cb.bvalid<=1'b0;
	@(vif.r_drv_cb);
	vif.r_drv_cb.bresp<=1'b0;

	/////////////////////read address channel//////////
	
	@(vif.r_drv_cb);
	vif.r_drv_cb.arready<=1'b1;
		@(vif.r_drv_cb);
		wait(vif.r_drv_cb.arvalid);
			@(vif.r_drv_cb);
			vif.r_drv_cb.arready<=1'b0;
			vif.r_drv_cb.araddr<=rtrans.araddr;
			vif.r_drv_cb.arprot<=rtrans.arprot;
	@(vif.r_drv_cb);

	//////////////read data or response //////////////////

		@(vif.r_drv_cb);
		vif.r_drv_cb.rvalid<=1'b1;
		@(vif.r_drv_cb);
		wait(vif.r_drv_cb.rready);
		@(vif.r_drv_cb);
		vif.r_drv_cb.rresp<=1'b1;

		vif.r_drv_cb.rdata<=rtrans.rdata;
		@(vif.r_drv_cb);


		num_sent1++;
		seq_item_port.item_done();
	end

end
endtask
*/
////////////////Repoprt Phase/////////////////////////////

function void report_phase(uvm_phase phase);
	   `uvm_info(get_type_name(), $sformatf("Report: FIFO RX DRIVER SENT %0d packets", num_sent1), UVM_LOW)
endfunction: report_phase

endclass  




